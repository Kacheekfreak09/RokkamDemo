�I�   } � eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffeefffffffffffeeeefeeeeeeeeeeeeeeeefeeeeeeeeeefeeeeeeeeffffffffffffgfffffffffffffffffffeefffeeeeeeeeeeeeeeeeeefeeeeeeeeeeeefeeeeffffffffffffffgggffffffffffffffffffeeffeeeeeeeeeeefffeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffgggggfffffgggggffffffffffeefeeeeeeeeeeeeeefffeeeeeeeeefeffeeeeeeeeeeeeffffffffffffffffffgNNNggggggggggggffffgffffeffeeeeeeeeeeeeeefffffeeeeeeefffffffeeeeeeeeeeeeeeeffffffffffefffgNNNNNggNNNNNNgggggggfgffeffeeeeeeeeeeeeeeeeeeefffffeeeeeeeffffffffffffeeeeeeeeeeeeeeeefggggffffffffggggNNNNNNNNNNgggggNNggffffeeefffeeeeeeeeeeeeeeeeeeeeffffeeeeeeefffffffffeeeffeeeeeeeeeeeefNNgggffffffffffgggNNNNNNNgggggNNNgggfffeeeffffeeeeeeeeeeeeeeeeeeeeeefffffeeeeeeeefffffffeeefffffffeeeeeeefNNNggffffffffffffggNNNNNNggggNNgggggfffeeeffffffeeeeeeeeeeeeeeeeeeeeeeefffffeeeeeeeeeffffffeeeeeffffeeeeeeeefgNNNggfffffffffffffggNNNNNggggNggggggffffeeefffffffeeeeeeeeeeeeeeeeeeeeeeeeefffffeeeeeeeeeeeffeeeeeffeeeeeeefggggggffffffeefffffffffgNNNNNNgffgggggggfffffeeeeefffffffeeeeeeeeeefeeffeeffeeeeeeeeeefffffeeeeeeeeeeeeeeeeeeeeeeeffffgggfffeeeeefffffffffggNNNNNggffffffffffffffffeeefffffffffeeeeeeeeeefffffeeeffeeeeeffffeeeefffffffeeeeeeeeeeeeeeeeeeeeeeeffffffggfeeeeeefffffffffggNNNNggffffffffffffffffffeffffffffffeeeeeeeeeefffffffeeeffeeeeeeffffffffffffffffeeeeeeeeeeeeefeeeeeeeefffffffffffffffffffffffffgggNgggffffffffeefffffffffffffffffffeeeeeeeefffffffffffffffeeeeeeeeffffffffffffffffeeeeeeeeeeefeeeefeeeeeffffffffffffffffeffffffffggggggffffffffeeeffffffffffffffffffeeeeeeeffffffffffffffeeefffeeeeeeefffffffffffffffffeeeeeeeeeeeeeeefffffffeeeffffffffffffffffffffffgggggfffffffffffffeefffgfffffffffffeeeeffffffffffffffffeeeeeeeeeefffffeeeeeeffffffgfffffffffffeeeeeeeeeeeeeeeeefffffeeeefffffffffffffffgggffffffffffffffffffffffffffggfffffffffeeeeffffffffffffffffffeeefeeeeeeefffffeeeeeffffggggfffffeefffeeeeeeeeeeeeeeeeeeeeefeeeeeeffffggfffffffffgggfffffffffffffffffffffffffffgffffffeeeeeeeffffffffffffffffffffffffffefffffffeeeeeefggggggfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffgggfffffffgggggffffffffffffffffffffffffffgffffffeeeeeeefffffffffffffffffffffffffffffffffffeeeeeffgNNNggffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffggggffffffgggggffffffffffggfffffffffeffffffffffeeeeeeeeeeeeefffffffffffffffffffffffffffffffeeeeffgNNNggfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffggfffffffffggfffffffffffggffffffffffffffffffffeeeeeeeeeeeeeffffffffffffffgffffffffffffffeeefffggNNggfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeffefffffffffMgffffffffffffffffffffggNggfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeefffeefffggffffffffffeeeeffffffgfgfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeefffffffffffffeeeeefffffgfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffefffeffffffffffeeffffffffffffffffffffffeeeeeeeeeeeeefffffffffffffffeeeeeffffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffeeeefffffffffffffffffffffeeeeeeeeeffffffffffffffffffeeefffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffeeeeeeefffffffeeeeeefffffeeeeeeeeeeeeefffffffffffffffeeefffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffeeeeeeeffffeeeeeeeeeeeeeffffeeeeffffeffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefeeeeeeeeeeefffeeeeeeeeeeeeeeeffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffeeeeeeeeeeeeeeeeffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffeeeeeeeeeeeeeefeeeeeeeeeeeeeeeeeeeeefffffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffeeeeeeffffeeeeeeeeeeeeeeeeeeeeeeeeeffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffeeeeeeeeeeeeeeeeeeeeeeeefffeeeeeeeeeeeeefffffeeeeeeeeefeeeeeeeeeeefffffeeeeeeeefeeefeeeefffeeeeeeeefeeeeeeeeefeeeeeeefeeeeeeeeeeeeeeeeeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffeeeeeeefffffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeffeeeeeeffffffffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefeeeeeeffffffffffffffeeeeeffffffeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffeefffffffffffeeeeeeeeeeeeeeeeeeeefeeeeeeeeeefeeeeeeeeffffffffffffgffffffffffffffffffeeeefeeeeeeeeeeeeeeeeefeeeeeeeeeeeefeeeeffffffffffffffgggffffffffffffffffffeefffeeeeeeffeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffgggggfffffgggggffffffeeffeeeeeeeeeeefffeeeeeeeeefeffeeeeeeeeeeeeffffffffffffffffffgNNNggggggggggggfffffffffeefeeeeeeeeeeeeeeffffeeeeeeefffffffeeeeeeeeeeeeeeeffffffffffefffgNNNNNggNNNNNNgggggggffffeffeeeeeeeeeeeeeefffffeeeeeeeffffffffffffeeeeeeeeeeeeeeeefggggffffffffggggNNNNNNNNNNggggggfgffeffeeeeeeeeeeeeeeeeeeefffffeeeeeeefffffffffeeeffeeeeeeeeeeeefNNgggffffffffffgggNNNNNNNgggggNNNggffffeeefffeeeeeeeeeeeeeeeeeeeefffffeeeeeeeefffffffeeefffffffeeeeeeefNNNggffffffffffffggNNNNNNggggNNNNgggfffeeeffffeeeeeeeeeeeeeeeeeeeeeefffffeeeeeeeeeffffffeeeeeffffeeeeeeeefgNNNggfffffffffffffggNNNNNggggNggggggfffeeeffffffeeeeeeeeeeeeeeeeeeeeeeefffffeeeeeeeeeeeffeeeeeffeeeeeeefggggggffffffeefffffffffgNNNNNNgffgggggggffffeeefffffffeeeeeeeeeeeeeeeeeeeeeeeeefffffeeeeeeeeeeeeeeeeeeeeeeeffffgggfffeeeeefffffffffggNNNNNggfffgggggfffffeeeeefffffffeeeeeeeeeefeeffeeffeeeeeeeeeeffffeeeeeeeeeeeeeeeeeeeeeeeffffffggfeeeeeefffffffffggNNNNggfffffffffffffffffeeefffffffffeeeeeeeeeefffffeeeffeeeeeffffeeeeffffffffeeeeeeeeeeeeefeeeeeeeefffffffffffffffffffffffffgggNgggffffffffffffffffffeffffffffffeeeeeeeeeefffffffeeeffeeeeeeffffffffffffffffeeeeeeeeeeefeeeefeeeeeffffffffffffffffeffffffffggggggfffffffffeefffffffffffffffffffeeeeeeeefffffffffffffffeeeeeeeeffffffffffffffffeeeeeeeeeeeeeeefffffffeeeffffffffffffffffffffffgggggffffffffeeeffffffffffffffffffeeeeeeeffffffffffffffeeefffeeeeeeefffffffffffffffffeeeeeeeeeeeeeeeeefffffeeeefffffffffffffffgggffffffffffffffffffffffeefffgfffffffffffeeeeffffffffffffffffeeeeeeeeeefffffeeeeeeffffffgfffffffefffeeeeeeeeeeeeeeeeeeeeefeeeeeeffffggfffffffffgggffffffffffffffffffffffffffggfffffffffeeeeffffffffffffffffffeeefeeeeeeefffffeeeeeffffggggfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffgggfffffffgggggffffffffffffffffffffffffffgffffffeeeeeeeffffffffffffffffffffffffffefffffffeeeeeefggggggfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffggggffffffgggggffffffffffggffffffffffffffgffffffeeeeeeefffffffffffffffffffffffffffffffffffeeeeeffgNNNggffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffggfffffffffggfffffffffffggfffffffffeffffffffffeeeeeeeeeeeeefffffffffffffffffffffffffffffffeeeeffgNNNggfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeffffffffffffffgffffffffffffffeeefffggNNggfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeffefffffffffMgffffffffffffffffffffggNggfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeefffeefffggffffffffffeeeeffffffgfgfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffefffeffffffffffeeffffffffffffffffffffffffeeeeeeeeeeeeeeeeeefffffffffffffeeeeefffffgfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffeeeefffffffffffffffffffffeeeeeeeeeeeeefffffffffffffffeeeeeffffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffeeeeeeeffffffffffffffffffffeeeeeeeeeffffffffffffffffffeeefffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffeeeeeeefffffeeeeeeeeeeeeefffffffffffffffeeefffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefeeeeeeeeeeffffeeeeeeeeeeeeeffffeeeeffffeffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffeeeeeeeeeeeeeeeffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffeeeeeeeeeeeeeeeeffeeeeeeeeeeeeeeeeeeeeefffeeeeeeeeeeeeeefeeeeeeeeeeeeeeeeeeefffffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeefffeeeeeeffffeeeeeeeeeeeeeeeeeeeeeeeeeffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffeeeeeeeeeeeeeeeeeeeeeeeeeefffeeeeeeeeeeefffffeeeeeeeeefeeeeeeeefffffeeeeeeeefeeefeeefffeeeeeeeefeeeeeeeeeeeeefeeeeeeefeeeeeeeeeeeeeeeeeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffeeeeeeefffffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeffeeeeeeffffffffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefeeeeeeffffffffffffffeeeeeffffffeef                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            